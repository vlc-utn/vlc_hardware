** Profile: "AC-AC"  [ e:\onedrive\universidad\utn\materias\6\proyecto_final\kicad\vlc_hardware\vlc_hardware\transmitter\fca\simulations\opa2675\lumicom_trans-pspicefiles\ac\ac.sim ] 

** Creating circuit file "AC.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Profile Libraries :
* Local Libraries :
* From [PSPICE NETLIST] section of C:\cds_spb_home\cdssetup\OrCAD_PSpiceTIPSpice_Install\23.1.0\PSpice.ini file:
.lib "nom_pspti.lib" 
.lib "nom.lib" 

*Analysis directives: 
.AC DEC 10 1k 10G
.OPTIONS ADVCONV
.OPTIONS FILEMODELSEARCH
.PROBE64 V(alias(*)) I(alias(*)) W(alias(*)) D(alias(*)) NOISE(alias(*)) 
.INC "..\AC.net" 


.END
