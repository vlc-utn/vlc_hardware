** Profile: "Noise-Noise"  [ E:\Onedrive\Universidad\UTN\Materias\6\proyecto_final\Simulaciones\PSpice\LMH34400\Archive\lmh34400-PSpiceFiles\Noise\Noise.sim ] 

** Creating circuit file "Noise.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Profile Libraries :
* Local Libraries :
.LIB "../../../LMH34400.lib" 
* From [PSPICE NETLIST] section of C:\cds_spb_home\cdssetup\OrCAD_PSpiceTIPSpice_Install\23.1.0\PSpice.ini file:
.lib "E:\Onedrive\Universidad\UTN\Materias\6\proyecto_final\Simulaciones\Modelos\Leds\Led_Chino.lib" 
.lib "nom_pspti.lib" 
.lib "nom.lib" 

*Analysis directives: 
.AC DEC 100 1K 10G
.NOISE V([OUT]) I_I1 1K
.OPTIONS ADVCONV
.OPTIONS FILEMODELSEARCH
.PROBE64 V(alias(*)) I(alias(*)) W(alias(*)) D(alias(*)) NOISE(alias(*)) 
.INC "..\Noise.net" 


.END
