** Profile: "AC-AC"  [ E:\Onedrive\Universidad\UTN\Materias\6\proyecto_final\Kicad\vlc_hardware\vlc_hardware\Transmitter\FCA\Simulations\OPA2675\lumicom_trans-pspicefiles\ac\ac.sim ] 

** Creating circuit file "AC.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Profile Libraries :
* Local Libraries :
.LIB "../../../library/infineon-rftransistor-spice.lib-sm-v02_10-en.lib" 
* From [PSPICE NETLIST] section of C:\cds_spb_home\cdssetup\OrCAD_PSpiceTIPSpice_Install\23.1.0\PSpice.ini file:
.lib "nom_pspti.lib" 
.lib "nom.lib" 

*Analysis directives: 
.AC DEC 100 1k 10G
.OPTIONS ADVCONV
.OPTIONS FILEMODELSEARCH
.PROBE64 V(alias(*)) I(alias(*)) W(alias(*)) D(alias(*)) NOISE(alias(*)) 
.INC "..\AC.net" 


.END
